library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Sparcv8Monocycle is
end Sparcv8Monocycle;

architecture Behavioral of Sparcv8Monocycle is

begin


end Behavioral;