library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity RF_Mux is
    Port ( RfDest : in  STD_LOGIC;
           RD : in  STD_LOGIC;
           nRD : out  STD_LOGIC_VECTOR (5 downto 0));
end RF_Mux;

architecture Behavioral of RF_Mux is

begin

process(RfDest, RD)
begin
	if (RfDest = '1') then
	end if;
end process;

end Behavioral;