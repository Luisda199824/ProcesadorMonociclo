library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity SignExtender is
    Port ( A : in  STD_LOGIC_VECTOR (12 downto 0);
           SEOut : out  STD_LOGIC_VECTOR (31 downto 0));
end SignExtender;

architecture Behavioral of SignExtender is

signal most : std_logic := '0'; -- Se�al que toma el bit m�s significativo de A
signal aux : std_logic_vector(31 downto 0) := (others => '0');

begin

most <= A(12);

process(A)
	begin
		if (most = '0') then
			SEOut <= "0000000000000000000"&A;
		else
			SEOut <= "1111111111111111111"&A;
		end if;
	end process;

end Behavioral;